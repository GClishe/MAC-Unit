`timescale 1ns/1ps

/*
 For this project, I will first store matrices written in A.mem and B.mem (potentially more later) to FPGA ROM.
 Then, upon a button press on the FPGA, matrices will be read and fed into 
*/
module matmul_top.sv(



);






endmodule 